// mfp_ahb_gpio.v
//
// General-purpose I/O module for Altera's DE2-115 and 
// Digilent's (Xilinx) Nexys4-DDR board
// License: Ram Bhattarai, Srijana Sapkota, Surya Ravikumar
//

/*Register MAPPING

`define H_7SEG_ENABLE_ADDR		(32'h1f700000)     //Physical address of Seven Segment Digit Enable Register
`define H_7SEG_UPPER_ADDR		(32'h1f700004)     //Physical address of Seven Segment UPPER Register
`define H_7SEG_LOWER_ADDR		(32'h1f700008)     //Physical address of Seven Segment LOWER Register
`define H_7SEG_DP_ADDR		    (32'h1f70000C)     //Physical address of Seven Segment Decimal Point register

//FOR SEVEN SEGMENT DISPLAY
Below numbers are generated by extracting 5:2 bits from the above Registers

`define H_7SEGEN_IONUM  		(4'h0)          //Using the same idea of GPIO's for MAPPING 5:2 bits 
`define H_7SEGUPPER_IONUM  		(4'h1)   
`define H_7SEGLOWER_IONUM  	    (4'h2)   
`define H_7SEGEDECIMAL_IONUM  	(4'h3)

*/ 


`include "mfp_ahb_const.vh"

module mfp_ahb_seven(
    input                        HCLK,
    input                        HRESETn,
    input      [  3          :0] HADDR,
    input      [  1          :0] HTRANS,
    input      [ 31          :0] HWDATA,
    input                        HWRITE,
    input                        HSEL,
    
    //Enable signal for 8 digits
    output [7:0] dispenout,
    
    //DP, CA, CB, CC, CC, CD, CE, CF
    output [7:0] dispout        
);

  reg  [7:0]  H7SEG_EN;                      //Seven segment enable register
  reg  [7:0]  H7SEG_DP;                      //Seven Segment Decimal points
  reg  [63:0] HSEG_DIGITS;        			// Seven segment Containing the upper and lower digit register
  
  reg  [3:0]  HADDR_d;
  reg         HWRITE_d;
  reg         HSEL_d;
  reg  [1:0]  HTRANS_d;
  
  wire        we;                               // write enable

  // delay HADDR, HWRITE, HSEL, and HTRANS to align with HWDATA for writing
  always @ (posedge HCLK) 
  begin
    HADDR_d  <= HADDR;
	HWRITE_d <= HWRITE;
	HSEL_d   <= HSEL;
	HTRANS_d <= HTRANS;
  end
  
  
  // overall write enable signal
  assign we = (HTRANS_d != `HTRANS_IDLE) & HSEL_d & HWRITE_d;

    always @(posedge HCLK or negedge HRESETn)
    begin
    
       if (~HRESETn)
            begin
                    H7SEG_EN <= 8'hff;
                    H7SEG_DP <= 8'hff;
                    HSEG_DIGITS<=64'hffffffff;
                
            end 
       else if (we)
         case (HADDR_d)
             //Based on the IOnumbers, select the hardware address
            `H_7SEGEN_IONUM        : H7SEG_EN    <= HWDATA[7:0];        
            `H_7SEGEDECIMAL_IONUM  : H7SEG_DP    <= HWDATA[7:0];
            `H_7SEGLOWER_IONUM     : HSEG_DIGITS[31:0] <= HWDATA; 
            `H_7SEGUPPER_IONUM     : HSEG_DIGITS[63:32] <= HWDATA;
            default:
            begin
                H7SEG_EN<= H7SEG_EN;
                HSEG_DIGITS<=HSEG_DIGITS;
                H7SEG_DP<=H7SEG_DP;  
            end
         endcase

    end
  
   
    //Instantiate the seven segment timer module
    mfp_ahb_sevensegtimer seven_segment_timer (.clk(HCLK), .resetn(HRESETn),.EN(H7SEG_EN),.DIGITS({HSEG_DIGITS}),
                                               .dp(H7SEG_DP),.DISPENOUT(dispenout),.DISPOUT(dispout));
endmodule

